
module unsaved (
	clk_clk,
	reset_reset_n,
	output_readra);	

	input		clk_clk;
	input		reset_reset_n;
	output		output_readra;
endmodule
